*** START IDEAL 10-BIT ADC Subcircuit ******************************
.subckt ADC10bit VDD VREFP VREFM Vin B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 CLOCK

* Set up common mode voltage
BCM VCM 0 V=(V(VREFP)-V(VREFM))/2

* Set up logic switching point
R3 VDD VTRIP 100MEG
R4 VTRIP 0 100MEG

* Ideal input sample and hold
XSH VDD VTRIP VIN OUTSH CLOCK SAMPHOLD

* Level shift by VREFM and 1/2LSB
BPIP PIPIN 0 V=V(OUTSH)-V(VREFM)+((V(VREFP)-V(VREFM))/2^11) ; 2^11 for 10-bit ADC

* 10-bit pipeline ADC
X9 VDD VTRIP VCM PIPIN B9 VOUT9 ADCBIT
X8 VDD VTRIP VCM VOUT9 B8 VOUT8 ADCBIT
X7 VDD VTRIP VCM VOUT8 B7 VOUT7 ADCBIT
X6 VDD VTRIP VCM VOUT7 B6 VOUT6 ADCBIT
X5 VDD VTRIP VCM VOUT6 B5 VOUT5 ADCBIT
X4 VDD VTRIP VCM VOUT5 B4 VOUT4 ADCBIT
X3 VDD VTRIP VCM VOUT4 B3 VOUT3 ADCBIT
X2 VDD VTRIP VCM VOUT3 B2 VOUT2 ADCBIT
X1 VDD VTRIP VCM VOUT2 B1 VOUT1 ADCBIT
X0 VDD VTRIP VCM VOUT1 B0 VOUT0 ADCBIT
.ends

* Ideal Sample and Hold subcircuit
.SUBCKT SAMPHOLD VDD VTRIP Vin Vout CLOCK
Ein Vinbuf 0 Vin Vinbuf 100MEG
S1 Vinbuf VinS VTRIP CLOCK switmod
Cs1 VinS 0 1e-10
S2 VinS Vout1 CLOCK VTRIP switmod
Cout1 Vout1 0 1e-16
Eout Vout 0 Vout1 0 1
.model switmod SW
.ends

* Pipeline stage
.SUBCKT ADCBIT VDD VTRIP VCM VIN BITOUT VOUT
S1 VDD BITOUT VIN VCM switmod
S2 0 BITOUT VCM VIN switmod
Eouth Vinh 0 VIN VCM 2
Eoutl Vinl 0 VIN 0 2
S3 Vinh VOUT BITOUT VTRIP switmod
S4 Vinl VOUT VTRIP BITOUT switmod
.model switmod SW
.ends

*** END ADC Subcircuit *************************************



*** Start Ideal 10-bit DAC Subcircuit *************************
.subckt DAC10bit VDD VREFP VREFM Vout B9 B8 B7 B6 B5 B4 B3 B2 B1 B0
*Generate Logic switching point, or trip, voltage
R1 VDD trip 100MEG
R2 trip 0 100MEG
*Change input logic signals into logic 0s or 1s
X9 trip B9 B9L Bitlogic
X8 trip B8 B8L Bitlogic
X7 trip B7 B7L Bitlogic
X6 trip B6 B6L Bitlogic
X5 trip B5 B5L Bitlogic
X4 trip B4 B4L Bitlogic
X3 trip B3 B3L Bitlogic
X2 trip B2 B2L Bitlogic
X1 trip B1 B1L Bitlogic
X0 trip B0 B0L Bitlogic
*Nonlinear dependent source, B, for generating the DAC output
Bout Vout 0 V=((v(vrefp)-v(vrefm))/1024)*(v(B9L)*512+v(B8L)*256+v(B7L)*128+v(B6L)*64+v(B5L)*32+v(B4L)*16+v(B3L)*8+v(B2L)*4+v(B1L)*2+v(B0L))+v(vrefm)
.ends
.subckt Bitlogic trip BX BXL
Vone one 0 DC 1
SH one BXL BX trip Switmod
SL 0 BXL trip BX Switmod
.model switmod SW
.ends
*** END DAC Subcircuit *************************************


*Simulation
X_myADC vdd vrefp vrefm vin b9 b8 b7 b6 b5 b4 b3 b2 b1 b0 clk ADC10bit

X_myDAC vdd vrefp vrefm vout b9 b8 b7 b6 b5 b4 b3 b2 b1 b0 DAC10bit

			  ; offset amp freq
V1 vin 0 DC 0 SIN(2.5 2.5 10653.40909)

V2 vdd 0 DC 5

V3 vrefp 0 DC 5

V4 vrefm 0 DC 0
; Vinit Von Tdelay Trise Tfall Ton Tperiod
V5 clk 0 pulse(0 5 0 1ns 1ns 0.55us 1.1us)

.tran 282.7us

